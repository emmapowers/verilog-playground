// config.svh
`ifndef CONFIG_SVH
`define CONFIG_SVH

`define CLOCK_FREQ_HZ 100_000_000  // 100 MHz
`define MS (`CLOCK_FREQ_HZ / 1000)  // Clock cycles in 1 Ms

`endif  // CONFIG_SVH
