package constants;

localparam int unsigned CLOCK_FREQ_HZ=100_000_000;  // 100 MHz
localparam int unsigned MS=(CLOCK_FREQ_HZ / 1000);  // Clock cycles in 1 Ms

endpackage